`timescale 1ns / 1ps

module tb_fan_adder_multi();
parameter DW_DATA = 8;
parameter DW_ROW = 4;
parameter DW_CTRL = 4;
parameter DW_LINE = DW_DATA + DW_ROW + DW_CTRL;
parameter NUM_IN = 2;

reg clk;
reg rst;
reg [NUM_IN*DW_LINE-1:0] in;
wire [NUM_IN*DW_LINE-1:0] out;

initial begin
    clk = 1'b1;
end
always #5 clk = ~clk;

initial begin
//    #10 // 111 110 
//    in = {16'b1010_0000_00000001, 16'b1000_0000_00000010, 167'b1000_0000_00000101, 16'b1000_0000_00010010, 16'b1001_0000_00100001, 16'b0100_0000_00000010};
//    #10 // 001 100
//    in = {16'b0100_00010_00000000, 16'b0000_0010_00100000, 16'b1000_0001_00000010, 16'b1001_0001_00000100, 16'b0100_0000_00000001, 16'b0000_0000_10000000};
    #10
    rst = 1'b1;
    in = 0;
    #10 // 11 10 add
    rst = 1'b0;
    // in = {16'b1010_0000_00000001, 16'b0000_0000_000000101, 16'b1001_0000_00100001, 16'b0111_0000_00000010};
    in = {16'b1010_0000_00000001, 16'b1001_0000_00000010};
    #30 // 01 10 bypass
    // in = {16'b0000_0010_00100000, 16'b1000_0010_00000010, 16'b1001_0001_00000100, 16'b0100_0000_00000001};
    in = {16'b1010_0001_00000001, 16'b1000_0001_00000010};
    #30
    // in = {16'b1010_0000_00000001, 16'b1000_0000_00000101, 16'b1001_0000_00100001, 16'b0100_0000_00000010};
    in = {16'b1010_0001_00000001, 16'b0111_0000_00000010};
//    #30
//    rst = 1'b0;
//    in = {16'b1010_0000_00000001, 16'b1001_0000_00000010};
//    #30
//    in = {16'b1010_0001_00000001, 16'b1000_0001_00000010};
    #100 $finish;
end

fan_adder_2to2 #(
    .DW_DATA(DW_DATA),
    .DW_ROW(DW_ROW),
    .DW_CTRL(DW_CTRL),
    .DW_LINE(DW_LINE)
) u_adder (
    .clk(clk),
//    .rst(rst),
    .in(in),
    .out(out)
);

endmodule   