`timescale 1ns / 1ps

module tb_ustc_fan();
parameter DW_DATA = 8;
parameter DW_ROW = 4;
parameter DW_CTRL = 4;
parameter DW_LINE = DW_DATA + DW_ROW + DW_CTRL;
//
parameter NUM_IN = 32;
parameter N_LEVELS = 5;

reg clk;
reg rst;
reg [NUM_IN*DW_LINE-1:0] in;
wire [NUM_IN*DW_LINE-1:0] out;

initial begin
    clk = 1'b1;
end
always #5 clk = ~clk;

initial begin
    in = 0;
    rst = 1'b1;
    #10
    rst = 1'b0;
    in = {16'b1010_0000_00011111, 16'b1000_0000_00011110, 16'b1001_0000_00011101,
          16'b1010_0001_00011100, 16'b1000_0001_00011011, 16'b1000_0001_00011010, 16'b1000_0001_00011001, 16'b1000_0001_00011000, 16'b1001_0001_00010111, 
          16'b1010_0010_00010110, 16'b1000_0010_00010101, 16'b1000_0010_00010100, 16'b1001_0010_00010011, 
          16'b1010_0011_00010010, 16'b1000_0011_00010001, 16'b1000_0011_00010000, 16'b1000_0011_00001111, 16'b1000_0011_00001110, 16'b1000_0011_00001101, 16'b1000_0011_00001100, 16'b1000_0011_00001011,
          16'b1000_0011_00001010, 16'b1000_0011_00001001, 16'b1001_0011_00001000,
          16'b1010_0100_00000111, 16'b1000_0100_00000110, 16'b1000_0100_00000101, 16'b1000_0100_00000100, 16'b1000_0100_00000011, 16'b1000_0100_00000010, 16'b1000_0100_00000001, 16'b1001_0100_00000000};
    #10 
    in = {16'b1010_0100_00000000, 16'b1000_0100_00000001, 16'b1000_0100_00000010, 16'b1000_0100_00000011, 16'b1000_0100_00000100, 16'b1000_0100_00000101, 16'b1000_0100_00000110, 16'b1001_0100_00000111,
          16'b1010_0011_00001000, 16'b1000_0011_00001001, 16'b1000_0011_00001010, 16'b1000_0011_00001011, 16'b1000_0011_00001100, 16'b1000_0011_00001101, 16'b1000_0011_00001110, 16'b1000_0011_00001111,
          16'b1000_0011_00010000, 16'b1000_0011_00010001, 16'b1001_0011_00010010, 
          16'b1010_0010_00010011, 16'b1000_0010_00010100, 16'b1000_0010_00010101, 16'b1001_0010_00010110, 
          16'b1010_0001_00010111, 16'b1000_0001_00011000, 16'b1000_0001_00011001, 16'b1000_0001_00011010, 16'b1000_0001_00011011, 16'b1001_0001_00011100, 
          16'b1010_0000_00011101, 16'b1000_0000_00011110, 16'b1001_0000_00011111};
    #10
    in = {16'b1010_0000_00011111, 16'b1000_0000_00011110, 16'b1001_0000_00011101,
          16'b1010_0001_00011100, 16'b1000_0001_00011011, 16'b1000_0001_00011010, 16'b1000_0001_00011001, 16'b1000_0001_00011000, 16'b1001_0001_00010111, 
          16'b1010_0010_00010110, 16'b1000_0010_00010101, 16'b1000_0010_00010100, 16'b1001_0010_00010011, 
          16'b1010_0011_00010010, 16'b1000_0011_00010001, 16'b1000_0011_00010000, 16'b1000_0011_00001111, 16'b1000_0011_00001110, 16'b1000_0011_00001101, 16'b1000_0011_00001100, 16'b1000_0011_00001011,
          16'b1000_0011_00001010, 16'b1000_0011_00001001, 16'b1001_0011_00001000,
          16'b1010_0100_00000111, 16'b1000_0100_00000110, 16'b1000_0100_00000101, 16'b1000_0100_00000100, 16'b1000_0100_00000011, 16'b1000_0100_00000010, 16'b1000_0100_00000001, 16'b1001_0100_00000000};
    #100 $finish;
end

ustc_fan #(
    .DW_DATA(DW_DATA),
    .DW_ROW(DW_ROW),
    .DW_CTRL(DW_CTRL),
    .DW_LINE(DW_LINE),
    .NUM_IN(NUM_IN)
) u_adder (
    .clk(clk),
    .rst(rst),
    .in(in),
    .out(out)
);

endmodule   